LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE symbols_7seg IS
	CONSTANT empty : STD_LOGIC_VECTOR(0 TO 6);
	
	CONSTANT H : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT L : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT O : STD_LOGIC_VECTOR(0 TO 6);
	
	CONSTANT zero : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT one : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT two : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT three : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT four : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT five : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT six : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT seven : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT eight : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT nine : STD_LOGIC_VECTOR(0 TO 6);

	CONSTANT A : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT B : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT C : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT D : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT E : STD_LOGIC_VECTOR(0 TO 6);
	CONSTANT F : STD_LOGIC_VECTOR(0 TO 6);
	
END PACKAGE symbols_7seg;

PACKAGE BODY symbols_7seg IS
	CONSTANT empty : STD_LOGIC_VECTOR(0 TO 6) := "1111111";

	CONSTANT H : STD_LOGIC_VECTOR(0 TO 6) := "1001000";
	CONSTANT L : STD_LOGIC_VECTOR(0 TO 6) := "1110001";
	CONSTANT O : STD_LOGIC_VECTOR(0 TO 6) := "0000001";
	
	CONSTANT zero : STD_LOGIC_VECTOR(0 TO 6) := "0000001";
	CONSTANT one : STD_LOGIC_VECTOR(0 TO 6) := "1001111";
	CONSTANT two : STD_LOGIC_VECTOR(0 TO 6) := "0010010";
	CONSTANT three : STD_LOGIC_VECTOR(0 TO 6) := "0000110";
	CONSTANT four : STD_LOGIC_VECTOR(0 TO 6) := "1001100";
	CONSTANT five : STD_LOGIC_VECTOR(0 TO 6) := "0100100";
	CONSTANT six : STD_LOGIC_VECTOR(0 TO 6) := "0100000";
	CONSTANT seven : STD_LOGIC_VECTOR(0 TO 6) := "0001111";
	CONSTANT eight : STD_LOGIC_VECTOR(0 TO 6) := "0000000";
	CONSTANT nine : STD_LOGIC_VECTOR(0 TO 6) := "0000100";
	
	CONSTANT A : STD_LOGIC_VECTOR(0 TO 6) := "0001000";
	CONSTANT B : STD_LOGIC_VECTOR(0 TO 6) := "1100000";
	CONSTANT C : STD_LOGIC_VECTOR(0 TO 6) := "0110001";
	CONSTANT D : STD_LOGIC_VECTOR(0 TO 6) := "1000010";
	CONSTANT E : STD_LOGIC_VECTOR(0 TO 6) := "0110000";
	CONSTANT F : STD_LOGIC_VECTOR(0 TO 6) := "0111000";
END PACKAGE BODY symbols_7seg;
